module MEM_WB(
input logic rst,
input logic clk,

input logic [4:0] RD_MEM_WB,
input logic REGFILE_WR_EN_MEM_WB,
input logic [31:0] REGFILE_IN_MEM_WB,

output logic [4:0] RD_REGFILE,
output logic REGFILE_WR_EN_REGFILE,
output logic [31:0] REGFILE_IN_REGFILE,
output logic [31:0] REGFILE_DATA_MEM_WB_REGISTER1,
output logic [31:0] REGFILE_DATA_MEM_WB_REGISTER2
);

logic [31:0] REGFILE_DATA_MEM_WB_REGISTER1_NEXT;
logic [31:0] REGFILE_DATA_MEM_WB_REGISTER2_NEXT;

always_comb begin
	RD_REGFILE = RD_MEM_WB;
	REGFILE_WR_EN_REGFILE = REGFILE_WR_EN_MEM_WB;
	REGFILE_IN_REGFILE = REGFILE_IN_MEM_WB;
if(REGFILE_WR_EN_REGFILE) begin
	REGFILE_DATA_MEM_WB_REGISTER1_NEXT = REGFILE_IN_MEM_WB;
	REGFILE_DATA_MEM_WB_REGISTER2_NEXT = REGFILE_DATA_MEM_WB_REGISTER1;
	end
else begin
		REGFILE_DATA_MEM_WB_REGISTER1_NEXT = REGFILE_DATA_MEM_WB_REGISTER1 ;
		REGFILE_DATA_MEM_WB_REGISTER2_NEXT = REGFILE_DATA_MEM_WB_REGISTER2 ;
	end
end

always_ff@(posedge clk)
begin

		REGFILE_DATA_MEM_WB_REGISTER1 <= REGFILE_DATA_MEM_WB_REGISTER1_NEXT ;
		REGFILE_DATA_MEM_WB_REGISTER2 <= REGFILE_DATA_MEM_WB_REGISTER2_NEXT ;

end

endmodule : MEM_WB